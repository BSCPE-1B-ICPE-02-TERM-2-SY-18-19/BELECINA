CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 7 120 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
176 80 1364 707
76546066 0
0
6 Title:
5 Name:
0
0
0
11
6 74112~
219 507 329 0 7 32
0 3 17 4 17 3 18 8
0
0 0 4704 0
5 74112
4 -60 39 -52
3 U6B
22 -61 43 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 10 11 13 12 14 7 9 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 2 5 0
1 U
6316 0 0
2
43528.9 10
0
6 74112~
219 368 329 0 7 32
0 3 16 4 16 3 19 5
0
0 0 4704 0
5 74112
4 -60 39 -52
3 U6A
22 -61 43 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 4 3 1 2 15 6 5 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 1 5 0
1 U
8734 0 0
2
43528.9 9
0
6 74112~
219 227 329 0 7 32
0 3 7 4 7 3 20 6
0
0 0 4704 0
5 74112
4 -60 39 -52
3 U4B
22 -61 43 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 10 11 13 12 14 7 9 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 2 4 0
1 U
7988 0 0
2
43528.9 8
0
6 74112~
219 123 328 0 7 32
0 3 3 4 3 3 21 7
0
0 0 4704 0
5 74112
4 -60 39 -52
3 U4A
22 -61 43 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 4 3 1 2 15 6 5 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 1 4 0
1 U
3217 0 0
2
43528.9 7
0
2 +V
167 123 215 0 1 3
0 3
0
0 0 54240 0
3 10V
-11 -22 10 -14
2 V2
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3965 0 0
2
43528.9 6
0
7 Ground~
168 686 118 0 1 3
0 2
0
0 0 53344 180
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
8239 0 0
2
43528.9 5
0
9 CC 7-Seg~
183 686 218 0 17 19
10 9 10 11 12 13 14 15 22 2
1 1 1 0 0 0 0 2
0
0 0 21104 0
5 REDCC
16 -41 51 -33
5 DISP1
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 1 0 0 0
4 DISP
828 0 0
2
43528.9 4
0
9 2-In AND~
219 296 195 0 3 22
0 7 6 16
0
0 0 608 0
6 74LS08
-21 -24 21 -16
3 U5A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 3 0
1 U
6187 0 0
2
43528.9 3
0
9 2-In AND~
219 432 204 0 3 22
0 16 5 17
0
0 0 608 0
6 74LS08
-21 -24 21 -16
3 U5B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 3 0
1 U
7107 0 0
2
43528.9 2
0
6 74LS48
188 593 411 0 14 29
0 8 5 6 7 23 24 15 14 13
12 11 10 9 25
0
0 0 4832 0
7 74LS248
-24 -60 25 -52
2 U3
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
119 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %14i]
+ [%16bo %1o %2o %3o %4o %5o %6o %14o %7o %8o %9o %10o %11o %12o %13o] %M
0
12 type:digital
5 DIP16
29

0 6 2 1 7 3 5 14 15 9
10 11 12 13 4 6 2 1 7 3
5 14 15 9 10 11 12 13 4 0
65 0 0 512 1 0 0 0
1 U
6433 0 0
2
43528.9 1
0
7 Pulser~
4 47 375 0 10 12
0 26 27 4 28 0 0 5 5 1
7
0
0 0 4640 0
0
2 V1
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
8559 0 0
2
43528.9 0
0
36
3 4 0 0 0 16 0 9 1 0 0 4
453 204
469 204
469 311
483 311
1 7 0 0 0 16 0 10 1 0 0 4
561 375
545 375
545 293
531 293
0 1 0 0 0 16 0 0 1 27 0 4
368 240
368 253
507 253
507 266
0 2 0 0 0 16 0 0 1 22 0 2
450 293
483 293
7 2 0 0 0 16 0 2 9 0 0 4
392 293
402 293
402 213
408 213
0 2 0 0 0 16 0 0 2 34 0 3
334 293
334 293
344 293
2 7 0 0 0 16 0 3 4 0 0 4
203 293
161 293
161 292
147 292
7 2 0 0 0 16 0 3 8 0 0 4
251 293
264 293
264 204
272 204
1 4 0 0 0 16 0 8 3 0 0 4
272 186
189 186
189 311
203 311
1 1 0 0 0 16 0 4 5 0 0 2
123 265
123 224
0 1 0 0 0 16 0 0 4 0 0 2
123 257
123 265
2 4 0 0 0 16 0 4 4 0 0 4
99 292
80 292
80 310
99 310
1 9 0 0 0 16 0 6 7 0 0 2
686 126
686 176
3 1 0 0 0 16 0 8 9 0 0 2
317 195
408 195
13 1 0 0 0 16 0 10 7 0 0 3
625 429
665 429
665 254
12 2 0 0 0 16 0 10 7 0 0 3
625 420
671 420
671 254
11 3 0 0 0 16 0 10 7 0 0 3
625 411
677 411
677 254
10 4 0 0 0 16 0 10 7 0 0 3
625 402
683 402
683 254
9 5 0 0 0 16 0 10 7 0 0 3
625 393
689 393
689 254
8 6 0 0 0 16 0 10 7 0 0 3
625 384
695 384
695 254
7 7 0 0 0 16 0 10 7 0 0 3
625 375
701 375
701 254
0 2 0 0 0 16 0 0 10 34 0 4
409 293
465 293
465 384
561 384
0 3 0 0 0 16 0 0 10 0 0 4
272 293
306 293
306 393
561 393
0 4 0 0 0 16 0 0 10 0 0 4
161 292
165 292
165 402
561 402
0 3 0 0 0 16 0 0 11 36 0 2
90 366
71 366
0 0 3 0 0 16 0 0 0 27 32 2
287 240
287 348
0 1 3 0 0 16 0 0 2 28 0 3
227 240
368 240
368 266
0 1 3 0 0 16 0 0 3 29 0 3
123 240
227 240
227 266
0 0 3 0 0 16 0 0 0 0 0 3
85 292
85 240
123 240
0 0 3 0 0 16 0 0 0 0 32 2
227 335
227 348
0 0 3 0 0 16 0 0 0 0 32 2
368 335
368 348
0 0 3 0 0 16 0 0 0 0 0 4
123 334
123 348
507 348
507 335
0 0 4 0 0 16 0 0 0 35 0 4
309 366
479 366
479 302
483 302
4 0 16 0 0 16 0 2 0 0 0 12
344 311
330 311
330 351
402 351
402 298
411 298
411 260
334 260
334 293
333 293
333 195
334 195
0 0 4 0 0 16 0 0 0 0 36 4
344 302
309 302
309 366
197 366
0 0 4 0 0 16 0 0 0 0 0 6
203 302
197 302
197 366
90 366
90 301
99 301
3
-35 0 0 0 400 0 0 0 0 3 2 1 82
7 Stencil
0 0 0 35
7 45 727 107
16 52 717 94
35 BINARY 4-BIT SYNCHRONOUS UP COUNTER
-21 0 0 0 700 255 0 0 0 3 2 1 2
17 SigismundoDiFanti
0 0 0 9
390 2 504 34
398 9 495 31
9 bscpe i-b
-21 0 0 0 700 255 0 0 0 3 2 1 2
17 SigismundoDiFanti
0 0 0 25
1 4 356 36
10 11 346 33
25 Ma. Jezabelle A. Belecina
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
